//////////////////////////////////////////////////////////////////////////////////
//
// This file is part of the N64 RGB/YPbPr DAC project.
//
// Copyright (C) 2015-2019 by Peter Bartmann <borti4938@gmx.de>
//
// N64 RGB/YPbPr DAC is free software: you can redistribute it and/or modify
// it under the terms of the GNU General Public License as published by
// the Free Software Foundation, either version 3 of the License, or
// any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program.  If not, see <http://www.gnu.org/licenses/>.
//
//////////////////////////////////////////////////////////////////////////////////
//
// Company:  Circuit-Board.de
// Engineer: borti4938
//
// Module Name:    font_rom
// Project Name:   N64 Advanced RGB/YPbPr DAC Mod
// Target Devices: Max10, Cyclone IV and Cyclone 10 LP devices
// Tool versions:  Altera Quartus Prime
// Description:    simple line-multiplying
//
// Features: ip independent implementation of font rom
//
// This file is auto generated by script/font2rom.m
//
//////////////////////////////////////////////////////////////////////////////////


module font_rom(
  CLK,
  nRST,
  char_addr,
  char_line,
  rden,
  rddata
);

input       CLK;
input       nRST;
input [6:0] char_addr;
input [3:0] char_line;
input       rden;

output reg [7:0] rddata;


reg [10:0] addr_r = 11'h00;
reg        rden_r =  1'b0;

always @(posedge CLK) begin
  addr_r <= {char_line,char_addr};
  rden_r <= rden;

  if (rden_r)
    case (addr_r)
      0000: rddata <= 000;
      0001: rddata <= 000;
      0002: rddata <= 000;
      0003: rddata <= 000;
      0004: rddata <= 000;
      0005: rddata <= 000;
      0006: rddata <= 000;
      0007: rddata <= 000;
      0008: rddata <= 000;
      0009: rddata <= 000;
      0010: rddata <= 000;
      0011: rddata <= 000;
      0012: rddata <= 000;
      0013: rddata <= 000;
      0014: rddata <= 000;
      0015: rddata <= 000;
      0016: rddata <= 000;
      0017: rddata <= 000;
      0018: rddata <= 000;
      0019: rddata <= 000;
      0020: rddata <= 000;
      0021: rddata <= 000;
      0022: rddata <= 000;
      0023: rddata <= 000;
      0024: rddata <= 000;
      0025: rddata <= 000;
      0026: rddata <= 000;
      0027: rddata <= 000;
      0028: rddata <= 000;
      0029: rddata <= 000;
      0030: rddata <= 000;
      0031: rddata <= 000;
      0032: rddata <= 000;
      0033: rddata <= 000;
      0034: rddata <= 000;
      0035: rddata <= 000;
      0036: rddata <= 012;
      0037: rddata <= 000;
      0038: rddata <= 000;
      0039: rddata <= 000;
      0040: rddata <= 000;
      0041: rddata <= 000;
      0042: rddata <= 000;
      0043: rddata <= 000;
      0044: rddata <= 000;
      0045: rddata <= 000;
      0046: rddata <= 000;
      0047: rddata <= 000;
      0048: rddata <= 000;
      0049: rddata <= 000;
      0050: rddata <= 000;
      0051: rddata <= 000;
      0052: rddata <= 000;
      0053: rddata <= 000;
      0054: rddata <= 000;
      0055: rddata <= 000;
      0056: rddata <= 000;
      0057: rddata <= 000;
      0058: rddata <= 000;
      0059: rddata <= 000;
      0060: rddata <= 000;
      0061: rddata <= 000;
      0062: rddata <= 000;
      0063: rddata <= 000;
      0064: rddata <= 000;
      0065: rddata <= 000;
      0066: rddata <= 000;
      0067: rddata <= 000;
      0068: rddata <= 000;
      0069: rddata <= 000;
      0070: rddata <= 000;
      0071: rddata <= 000;
      0072: rddata <= 000;
      0073: rddata <= 000;
      0074: rddata <= 000;
      0075: rddata <= 000;
      0076: rddata <= 000;
      0077: rddata <= 000;
      0078: rddata <= 000;
      0079: rddata <= 000;
      0080: rddata <= 000;
      0081: rddata <= 000;
      0082: rddata <= 000;
      0083: rddata <= 000;
      0084: rddata <= 000;
      0085: rddata <= 000;
      0086: rddata <= 000;
      0087: rddata <= 000;
      0088: rddata <= 000;
      0089: rddata <= 000;
      0090: rddata <= 000;
      0091: rddata <= 000;
      0092: rddata <= 000;
      0093: rddata <= 000;
      0094: rddata <= 008;
      0095: rddata <= 000;
      0096: rddata <= 012;
      0097: rddata <= 000;
      0098: rddata <= 000;
      0099: rddata <= 000;
      0100: rddata <= 000;
      0101: rddata <= 000;
      0102: rddata <= 000;
      0103: rddata <= 000;
      0104: rddata <= 000;
      0105: rddata <= 000;
      0106: rddata <= 000;
      0107: rddata <= 000;
      0108: rddata <= 000;
      0109: rddata <= 000;
      0110: rddata <= 000;
      0111: rddata <= 000;
      0112: rddata <= 000;
      0113: rddata <= 000;
      0114: rddata <= 000;
      0115: rddata <= 000;
      0116: rddata <= 000;
      0117: rddata <= 000;
      0118: rddata <= 000;
      0119: rddata <= 000;
      0120: rddata <= 000;
      0121: rddata <= 000;
      0122: rddata <= 000;
      0123: rddata <= 000;
      0124: rddata <= 000;
      0125: rddata <= 000;
      0126: rddata <= 000;
      0127: rddata <= 000;
      0128: rddata <= 000;
      0129: rddata <= 000;
      0130: rddata <= 126;
      0131: rddata <= 000;
      0132: rddata <= 008;
      0133: rddata <= 024;
      0134: rddata <= 024;
      0135: rddata <= 000;
      0136: rddata <= 000;
      0137: rddata <= 028;
      0138: rddata <= 028;
      0139: rddata <= 124;
      0140: rddata <= 060;
      0141: rddata <= 000;
      0142: rddata <= 254;
      0143: rddata <= 000;
      0144: rddata <= 064;
      0145: rddata <= 001;
      0146: rddata <= 024;
      0147: rddata <= 102;
      0148: rddata <= 254;
      0149: rddata <= 126;
      0150: rddata <= 000;
      0151: rddata <= 024;
      0152: rddata <= 024;
      0153: rddata <= 024;
      0154: rddata <= 000;
      0155: rddata <= 000;
      0156: rddata <= 000;
      0157: rddata <= 000;
      0158: rddata <= 000;
      0159: rddata <= 000;
      0160: rddata <= 000;
      0161: rddata <= 012;
      0162: rddata <= 102;
      0163: rddata <= 054;
      0164: rddata <= 012;
      0165: rddata <= 000;
      0166: rddata <= 014;
      0167: rddata <= 012;
      0168: rddata <= 048;
      0169: rddata <= 006;
      0170: rddata <= 000;
      0171: rddata <= 000;
      0172: rddata <= 000;
      0173: rddata <= 000;
      0174: rddata <= 000;
      0175: rddata <= 000;
      0176: rddata <= 062;
      0177: rddata <= 008;
      0178: rddata <= 030;
      0179: rddata <= 030;
      0180: rddata <= 048;
      0181: rddata <= 063;
      0182: rddata <= 028;
      0183: rddata <= 127;
      0184: rddata <= 030;
      0185: rddata <= 030;
      0186: rddata <= 000;
      0187: rddata <= 000;
      0188: rddata <= 048;
      0189: rddata <= 000;
      0190: rddata <= 006;
      0191: rddata <= 030;
      0192: rddata <= 062;
      0193: rddata <= 012;
      0194: rddata <= 063;
      0195: rddata <= 060;
      0196: rddata <= 031;
      0197: rddata <= 127;
      0198: rddata <= 127;
      0199: rddata <= 060;
      0200: rddata <= 051;
      0201: rddata <= 030;
      0202: rddata <= 120;
      0203: rddata <= 103;
      0204: rddata <= 015;
      0205: rddata <= 099;
      0206: rddata <= 099;
      0207: rddata <= 028;
      0208: rddata <= 063;
      0209: rddata <= 028;
      0210: rddata <= 063;
      0211: rddata <= 030;
      0212: rddata <= 063;
      0213: rddata <= 051;
      0214: rddata <= 051;
      0215: rddata <= 099;
      0216: rddata <= 051;
      0217: rddata <= 051;
      0218: rddata <= 127;
      0219: rddata <= 060;
      0220: rddata <= 000;
      0221: rddata <= 060;
      0222: rddata <= 028;
      0223: rddata <= 000;
      0224: rddata <= 012;
      0225: rddata <= 000;
      0226: rddata <= 007;
      0227: rddata <= 000;
      0228: rddata <= 056;
      0229: rddata <= 000;
      0230: rddata <= 028;
      0231: rddata <= 000;
      0232: rddata <= 007;
      0233: rddata <= 024;
      0234: rddata <= 048;
      0235: rddata <= 007;
      0236: rddata <= 030;
      0237: rddata <= 000;
      0238: rddata <= 000;
      0239: rddata <= 000;
      0240: rddata <= 000;
      0241: rddata <= 000;
      0242: rddata <= 000;
      0243: rddata <= 000;
      0244: rddata <= 000;
      0245: rddata <= 000;
      0246: rddata <= 000;
      0247: rddata <= 000;
      0248: rddata <= 000;
      0249: rddata <= 000;
      0250: rddata <= 000;
      0251: rddata <= 056;
      0252: rddata <= 024;
      0253: rddata <= 007;
      0254: rddata <= 206;
      0255: rddata <= 000;
      0256: rddata <= 000;
      0257: rddata <= 000;
      0258: rddata <= 195;
      0259: rddata <= 034;
      0260: rddata <= 028;
      0261: rddata <= 060;
      0262: rddata <= 060;
      0263: rddata <= 255;
      0264: rddata <= 255;
      0265: rddata <= 034;
      0266: rddata <= 034;
      0267: rddata <= 112;
      0268: rddata <= 102;
      0269: rddata <= 000;
      0270: rddata <= 198;
      0271: rddata <= 024;
      0272: rddata <= 096;
      0273: rddata <= 003;
      0274: rddata <= 060;
      0275: rddata <= 102;
      0276: rddata <= 219;
      0277: rddata <= 198;
      0278: rddata <= 000;
      0279: rddata <= 060;
      0280: rddata <= 060;
      0281: rddata <= 024;
      0282: rddata <= 000;
      0283: rddata <= 000;
      0284: rddata <= 000;
      0285: rddata <= 000;
      0286: rddata <= 008;
      0287: rddata <= 127;
      0288: rddata <= 000;
      0289: rddata <= 030;
      0290: rddata <= 102;
      0291: rddata <= 054;
      0292: rddata <= 062;
      0293: rddata <= 000;
      0294: rddata <= 027;
      0295: rddata <= 012;
      0296: rddata <= 024;
      0297: rddata <= 012;
      0298: rddata <= 000;
      0299: rddata <= 000;
      0300: rddata <= 000;
      0301: rddata <= 000;
      0302: rddata <= 000;
      0303: rddata <= 064;
      0304: rddata <= 099;
      0305: rddata <= 012;
      0306: rddata <= 051;
      0307: rddata <= 051;
      0308: rddata <= 056;
      0309: rddata <= 003;
      0310: rddata <= 006;
      0311: rddata <= 099;
      0312: rddata <= 051;
      0313: rddata <= 051;
      0314: rddata <= 000;
      0315: rddata <= 000;
      0316: rddata <= 024;
      0317: rddata <= 000;
      0318: rddata <= 012;
      0319: rddata <= 051;
      0320: rddata <= 099;
      0321: rddata <= 030;
      0322: rddata <= 102;
      0323: rddata <= 102;
      0324: rddata <= 054;
      0325: rddata <= 070;
      0326: rddata <= 102;
      0327: rddata <= 102;
      0328: rddata <= 051;
      0329: rddata <= 012;
      0330: rddata <= 048;
      0331: rddata <= 102;
      0332: rddata <= 006;
      0333: rddata <= 119;
      0334: rddata <= 099;
      0335: rddata <= 054;
      0336: rddata <= 102;
      0337: rddata <= 054;
      0338: rddata <= 102;
      0339: rddata <= 051;
      0340: rddata <= 045;
      0341: rddata <= 051;
      0342: rddata <= 051;
      0343: rddata <= 099;
      0344: rddata <= 051;
      0345: rddata <= 051;
      0346: rddata <= 115;
      0347: rddata <= 012;
      0348: rddata <= 001;
      0349: rddata <= 048;
      0350: rddata <= 054;
      0351: rddata <= 000;
      0352: rddata <= 024;
      0353: rddata <= 000;
      0354: rddata <= 006;
      0355: rddata <= 000;
      0356: rddata <= 048;
      0357: rddata <= 000;
      0358: rddata <= 054;
      0359: rddata <= 000;
      0360: rddata <= 006;
      0361: rddata <= 024;
      0362: rddata <= 048;
      0363: rddata <= 006;
      0364: rddata <= 024;
      0365: rddata <= 000;
      0366: rddata <= 000;
      0367: rddata <= 000;
      0368: rddata <= 000;
      0369: rddata <= 000;
      0370: rddata <= 000;
      0371: rddata <= 000;
      0372: rddata <= 004;
      0373: rddata <= 000;
      0374: rddata <= 000;
      0375: rddata <= 000;
      0376: rddata <= 000;
      0377: rddata <= 000;
      0378: rddata <= 000;
      0379: rddata <= 012;
      0380: rddata <= 024;
      0381: rddata <= 012;
      0382: rddata <= 091;
      0383: rddata <= 000;
      0384: rddata <= 000;
      0385: rddata <= 000;
      0386: rddata <= 129;
      0387: rddata <= 119;
      0388: rddata <= 062;
      0389: rddata <= 060;
      0390: rddata <= 126;
      0391: rddata <= 000;
      0392: rddata <= 000;
      0393: rddata <= 093;
      0394: rddata <= 093;
      0395: rddata <= 092;
      0396: rddata <= 102;
      0397: rddata <= 000;
      0398: rddata <= 254;
      0399: rddata <= 219;
      0400: rddata <= 112;
      0401: rddata <= 007;
      0402: rddata <= 126;
      0403: rddata <= 102;
      0404: rddata <= 219;
      0405: rddata <= 012;
      0406: rddata <= 000;
      0407: rddata <= 126;
      0408: rddata <= 126;
      0409: rddata <= 024;
      0410: rddata <= 012;
      0411: rddata <= 024;
      0412: rddata <= 000;
      0413: rddata <= 036;
      0414: rddata <= 008;
      0415: rddata <= 127;
      0416: rddata <= 000;
      0417: rddata <= 030;
      0418: rddata <= 102;
      0419: rddata <= 127;
      0420: rddata <= 003;
      0421: rddata <= 035;
      0422: rddata <= 027;
      0423: rddata <= 012;
      0424: rddata <= 012;
      0425: rddata <= 024;
      0426: rddata <= 102;
      0427: rddata <= 024;
      0428: rddata <= 000;
      0429: rddata <= 000;
      0430: rddata <= 000;
      0431: rddata <= 096;
      0432: rddata <= 115;
      0433: rddata <= 015;
      0434: rddata <= 051;
      0435: rddata <= 048;
      0436: rddata <= 060;
      0437: rddata <= 003;
      0438: rddata <= 003;
      0439: rddata <= 099;
      0440: rddata <= 051;
      0441: rddata <= 051;
      0442: rddata <= 028;
      0443: rddata <= 028;
      0444: rddata <= 012;
      0445: rddata <= 000;
      0446: rddata <= 024;
      0447: rddata <= 048;
      0448: rddata <= 099;
      0449: rddata <= 051;
      0450: rddata <= 102;
      0451: rddata <= 099;
      0452: rddata <= 102;
      0453: rddata <= 006;
      0454: rddata <= 070;
      0455: rddata <= 099;
      0456: rddata <= 051;
      0457: rddata <= 012;
      0458: rddata <= 048;
      0459: rddata <= 054;
      0460: rddata <= 006;
      0461: rddata <= 127;
      0462: rddata <= 103;
      0463: rddata <= 099;
      0464: rddata <= 102;
      0465: rddata <= 099;
      0466: rddata <= 102;
      0467: rddata <= 051;
      0468: rddata <= 012;
      0469: rddata <= 051;
      0470: rddata <= 051;
      0471: rddata <= 099;
      0472: rddata <= 051;
      0473: rddata <= 051;
      0474: rddata <= 025;
      0475: rddata <= 012;
      0476: rddata <= 003;
      0477: rddata <= 048;
      0478: rddata <= 099;
      0479: rddata <= 000;
      0480: rddata <= 000;
      0481: rddata <= 000;
      0482: rddata <= 006;
      0483: rddata <= 000;
      0484: rddata <= 048;
      0485: rddata <= 000;
      0486: rddata <= 006;
      0487: rddata <= 000;
      0488: rddata <= 006;
      0489: rddata <= 000;
      0490: rddata <= 000;
      0491: rddata <= 006;
      0492: rddata <= 024;
      0493: rddata <= 000;
      0494: rddata <= 000;
      0495: rddata <= 000;
      0496: rddata <= 000;
      0497: rddata <= 000;
      0498: rddata <= 000;
      0499: rddata <= 000;
      0500: rddata <= 006;
      0501: rddata <= 000;
      0502: rddata <= 000;
      0503: rddata <= 000;
      0504: rddata <= 000;
      0505: rddata <= 000;
      0506: rddata <= 000;
      0507: rddata <= 012;
      0508: rddata <= 024;
      0509: rddata <= 012;
      0510: rddata <= 115;
      0511: rddata <= 008;
      0512: rddata <= 000;
      0513: rddata <= 000;
      0514: rddata <= 165;
      0515: rddata <= 127;
      0516: rddata <= 127;
      0517: rddata <= 255;
      0518: rddata <= 255;
      0519: rddata <= 000;
      0520: rddata <= 255;
      0521: rddata <= 085;
      0522: rddata <= 069;
      0523: rddata <= 078;
      0524: rddata <= 102;
      0525: rddata <= 000;
      0526: rddata <= 198;
      0527: rddata <= 126;
      0528: rddata <= 124;
      0529: rddata <= 031;
      0530: rddata <= 024;
      0531: rddata <= 102;
      0532: rddata <= 219;
      0533: rddata <= 060;
      0534: rddata <= 000;
      0535: rddata <= 024;
      0536: rddata <= 024;
      0537: rddata <= 024;
      0538: rddata <= 006;
      0539: rddata <= 048;
      0540: rddata <= 003;
      0541: rddata <= 102;
      0542: rddata <= 028;
      0543: rddata <= 062;
      0544: rddata <= 000;
      0545: rddata <= 030;
      0546: rddata <= 036;
      0547: rddata <= 054;
      0548: rddata <= 003;
      0549: rddata <= 051;
      0550: rddata <= 014;
      0551: rddata <= 006;
      0552: rddata <= 006;
      0553: rddata <= 048;
      0554: rddata <= 060;
      0555: rddata <= 024;
      0556: rddata <= 000;
      0557: rddata <= 000;
      0558: rddata <= 000;
      0559: rddata <= 048;
      0560: rddata <= 123;
      0561: rddata <= 012;
      0562: rddata <= 048;
      0563: rddata <= 048;
      0564: rddata <= 054;
      0565: rddata <= 003;
      0566: rddata <= 003;
      0567: rddata <= 096;
      0568: rddata <= 051;
      0569: rddata <= 051;
      0570: rddata <= 028;
      0571: rddata <= 028;
      0572: rddata <= 006;
      0573: rddata <= 126;
      0574: rddata <= 048;
      0575: rddata <= 024;
      0576: rddata <= 123;
      0577: rddata <= 051;
      0578: rddata <= 102;
      0579: rddata <= 003;
      0580: rddata <= 102;
      0581: rddata <= 038;
      0582: rddata <= 038;
      0583: rddata <= 003;
      0584: rddata <= 051;
      0585: rddata <= 012;
      0586: rddata <= 048;
      0587: rddata <= 054;
      0588: rddata <= 006;
      0589: rddata <= 127;
      0590: rddata <= 111;
      0591: rddata <= 099;
      0592: rddata <= 102;
      0593: rddata <= 099;
      0594: rddata <= 102;
      0595: rddata <= 003;
      0596: rddata <= 012;
      0597: rddata <= 051;
      0598: rddata <= 051;
      0599: rddata <= 099;
      0600: rddata <= 030;
      0601: rddata <= 051;
      0602: rddata <= 024;
      0603: rddata <= 012;
      0604: rddata <= 006;
      0605: rddata <= 048;
      0606: rddata <= 000;
      0607: rddata <= 000;
      0608: rddata <= 000;
      0609: rddata <= 030;
      0610: rddata <= 062;
      0611: rddata <= 030;
      0612: rddata <= 062;
      0613: rddata <= 030;
      0614: rddata <= 006;
      0615: rddata <= 110;
      0616: rddata <= 054;
      0617: rddata <= 030;
      0618: rddata <= 060;
      0619: rddata <= 102;
      0620: rddata <= 024;
      0621: rddata <= 063;
      0622: rddata <= 031;
      0623: rddata <= 030;
      0624: rddata <= 059;
      0625: rddata <= 110;
      0626: rddata <= 055;
      0627: rddata <= 030;
      0628: rddata <= 063;
      0629: rddata <= 051;
      0630: rddata <= 051;
      0631: rddata <= 099;
      0632: rddata <= 099;
      0633: rddata <= 102;
      0634: rddata <= 063;
      0635: rddata <= 006;
      0636: rddata <= 024;
      0637: rddata <= 024;
      0638: rddata <= 000;
      0639: rddata <= 028;
      0640: rddata <= 000;
      0641: rddata <= 000;
      0642: rddata <= 129;
      0643: rddata <= 127;
      0644: rddata <= 127;
      0645: rddata <= 231;
      0646: rddata <= 255;
      0647: rddata <= 000;
      0648: rddata <= 000;
      0649: rddata <= 093;
      0650: rddata <= 069;
      0651: rddata <= 031;
      0652: rddata <= 060;
      0653: rddata <= 000;
      0654: rddata <= 198;
      0655: rddata <= 231;
      0656: rddata <= 127;
      0657: rddata <= 127;
      0658: rddata <= 024;
      0659: rddata <= 102;
      0660: rddata <= 222;
      0661: rddata <= 102;
      0662: rddata <= 000;
      0663: rddata <= 024;
      0664: rddata <= 024;
      0665: rddata <= 024;
      0666: rddata <= 127;
      0667: rddata <= 127;
      0668: rddata <= 003;
      0669: rddata <= 255;
      0670: rddata <= 028;
      0671: rddata <= 062;
      0672: rddata <= 000;
      0673: rddata <= 012;
      0674: rddata <= 000;
      0675: rddata <= 054;
      0676: rddata <= 030;
      0677: rddata <= 024;
      0678: rddata <= 095;
      0679: rddata <= 000;
      0680: rddata <= 006;
      0681: rddata <= 048;
      0682: rddata <= 255;
      0683: rddata <= 126;
      0684: rddata <= 000;
      0685: rddata <= 127;
      0686: rddata <= 000;
      0687: rddata <= 024;
      0688: rddata <= 107;
      0689: rddata <= 012;
      0690: rddata <= 024;
      0691: rddata <= 028;
      0692: rddata <= 051;
      0693: rddata <= 031;
      0694: rddata <= 031;
      0695: rddata <= 048;
      0696: rddata <= 030;
      0697: rddata <= 062;
      0698: rddata <= 000;
      0699: rddata <= 000;
      0700: rddata <= 003;
      0701: rddata <= 000;
      0702: rddata <= 096;
      0703: rddata <= 012;
      0704: rddata <= 123;
      0705: rddata <= 051;
      0706: rddata <= 062;
      0707: rddata <= 003;
      0708: rddata <= 102;
      0709: rddata <= 062;
      0710: rddata <= 062;
      0711: rddata <= 003;
      0712: rddata <= 063;
      0713: rddata <= 012;
      0714: rddata <= 048;
      0715: rddata <= 030;
      0716: rddata <= 006;
      0717: rddata <= 107;
      0718: rddata <= 127;
      0719: rddata <= 099;
      0720: rddata <= 062;
      0721: rddata <= 099;
      0722: rddata <= 062;
      0723: rddata <= 014;
      0724: rddata <= 012;
      0725: rddata <= 051;
      0726: rddata <= 051;
      0727: rddata <= 107;
      0728: rddata <= 012;
      0729: rddata <= 030;
      0730: rddata <= 012;
      0731: rddata <= 012;
      0732: rddata <= 012;
      0733: rddata <= 048;
      0734: rddata <= 000;
      0735: rddata <= 000;
      0736: rddata <= 000;
      0737: rddata <= 048;
      0738: rddata <= 102;
      0739: rddata <= 051;
      0740: rddata <= 051;
      0741: rddata <= 051;
      0742: rddata <= 031;
      0743: rddata <= 051;
      0744: rddata <= 110;
      0745: rddata <= 024;
      0746: rddata <= 048;
      0747: rddata <= 054;
      0748: rddata <= 024;
      0749: rddata <= 107;
      0750: rddata <= 051;
      0751: rddata <= 051;
      0752: rddata <= 102;
      0753: rddata <= 051;
      0754: rddata <= 118;
      0755: rddata <= 051;
      0756: rddata <= 006;
      0757: rddata <= 051;
      0758: rddata <= 051;
      0759: rddata <= 099;
      0760: rddata <= 054;
      0761: rddata <= 102;
      0762: rddata <= 049;
      0763: rddata <= 003;
      0764: rddata <= 000;
      0765: rddata <= 048;
      0766: rddata <= 000;
      0767: rddata <= 054;
      0768: rddata <= 000;
      0769: rddata <= 000;
      0770: rddata <= 189;
      0771: rddata <= 127;
      0772: rddata <= 062;
      0773: rddata <= 231;
      0774: rddata <= 126;
      0775: rddata <= 000;
      0776: rddata <= 000;
      0777: rddata <= 077;
      0778: rddata <= 069;
      0779: rddata <= 051;
      0780: rddata <= 024;
      0781: rddata <= 000;
      0782: rddata <= 198;
      0783: rddata <= 231;
      0784: rddata <= 124;
      0785: rddata <= 031;
      0786: rddata <= 024;
      0787: rddata <= 000;
      0788: rddata <= 216;
      0789: rddata <= 102;
      0790: rddata <= 000;
      0791: rddata <= 024;
      0792: rddata <= 024;
      0793: rddata <= 024;
      0794: rddata <= 006;
      0795: rddata <= 048;
      0796: rddata <= 003;
      0797: rddata <= 102;
      0798: rddata <= 062;
      0799: rddata <= 028;
      0800: rddata <= 000;
      0801: rddata <= 012;
      0802: rddata <= 000;
      0803: rddata <= 054;
      0804: rddata <= 048;
      0805: rddata <= 012;
      0806: rddata <= 123;
      0807: rddata <= 000;
      0808: rddata <= 006;
      0809: rddata <= 048;
      0810: rddata <= 060;
      0811: rddata <= 024;
      0812: rddata <= 000;
      0813: rddata <= 000;
      0814: rddata <= 000;
      0815: rddata <= 012;
      0816: rddata <= 111;
      0817: rddata <= 012;
      0818: rddata <= 012;
      0819: rddata <= 048;
      0820: rddata <= 127;
      0821: rddata <= 048;
      0822: rddata <= 051;
      0823: rddata <= 024;
      0824: rddata <= 051;
      0825: rddata <= 024;
      0826: rddata <= 000;
      0827: rddata <= 000;
      0828: rddata <= 006;
      0829: rddata <= 126;
      0830: rddata <= 048;
      0831: rddata <= 012;
      0832: rddata <= 123;
      0833: rddata <= 063;
      0834: rddata <= 102;
      0835: rddata <= 003;
      0836: rddata <= 102;
      0837: rddata <= 038;
      0838: rddata <= 038;
      0839: rddata <= 115;
      0840: rddata <= 051;
      0841: rddata <= 012;
      0842: rddata <= 051;
      0843: rddata <= 054;
      0844: rddata <= 070;
      0845: rddata <= 099;
      0846: rddata <= 123;
      0847: rddata <= 099;
      0848: rddata <= 006;
      0849: rddata <= 115;
      0850: rddata <= 054;
      0851: rddata <= 024;
      0852: rddata <= 012;
      0853: rddata <= 051;
      0854: rddata <= 051;
      0855: rddata <= 107;
      0856: rddata <= 030;
      0857: rddata <= 012;
      0858: rddata <= 006;
      0859: rddata <= 012;
      0860: rddata <= 024;
      0861: rddata <= 048;
      0862: rddata <= 000;
      0863: rddata <= 000;
      0864: rddata <= 000;
      0865: rddata <= 062;
      0866: rddata <= 102;
      0867: rddata <= 003;
      0868: rddata <= 051;
      0869: rddata <= 063;
      0870: rddata <= 006;
      0871: rddata <= 051;
      0872: rddata <= 102;
      0873: rddata <= 024;
      0874: rddata <= 048;
      0875: rddata <= 030;
      0876: rddata <= 024;
      0877: rddata <= 107;
      0878: rddata <= 051;
      0879: rddata <= 051;
      0880: rddata <= 102;
      0881: rddata <= 051;
      0882: rddata <= 110;
      0883: rddata <= 006;
      0884: rddata <= 006;
      0885: rddata <= 051;
      0886: rddata <= 051;
      0887: rddata <= 107;
      0888: rddata <= 028;
      0889: rddata <= 102;
      0890: rddata <= 024;
      0891: rddata <= 006;
      0892: rddata <= 024;
      0893: rddata <= 024;
      0894: rddata <= 000;
      0895: rddata <= 099;
      0896: rddata <= 000;
      0897: rddata <= 000;
      0898: rddata <= 153;
      0899: rddata <= 062;
      0900: rddata <= 028;
      0901: rddata <= 024;
      0902: rddata <= 024;
      0903: rddata <= 000;
      0904: rddata <= 000;
      0905: rddata <= 085;
      0906: rddata <= 093;
      0907: rddata <= 051;
      0908: rddata <= 126;
      0909: rddata <= 000;
      0910: rddata <= 230;
      0911: rddata <= 126;
      0912: rddata <= 112;
      0913: rddata <= 007;
      0914: rddata <= 126;
      0915: rddata <= 000;
      0916: rddata <= 216;
      0917: rddata <= 060;
      0918: rddata <= 127;
      0919: rddata <= 126;
      0920: rddata <= 024;
      0921: rddata <= 126;
      0922: rddata <= 012;
      0923: rddata <= 024;
      0924: rddata <= 127;
      0925: rddata <= 036;
      0926: rddata <= 062;
      0927: rddata <= 028;
      0928: rddata <= 000;
      0929: rddata <= 000;
      0930: rddata <= 000;
      0931: rddata <= 127;
      0932: rddata <= 048;
      0933: rddata <= 006;
      0934: rddata <= 051;
      0935: rddata <= 000;
      0936: rddata <= 012;
      0937: rddata <= 024;
      0938: rddata <= 102;
      0939: rddata <= 024;
      0940: rddata <= 000;
      0941: rddata <= 000;
      0942: rddata <= 000;
      0943: rddata <= 006;
      0944: rddata <= 103;
      0945: rddata <= 012;
      0946: rddata <= 006;
      0947: rddata <= 048;
      0948: rddata <= 048;
      0949: rddata <= 048;
      0950: rddata <= 051;
      0951: rddata <= 012;
      0952: rddata <= 051;
      0953: rddata <= 024;
      0954: rddata <= 028;
      0955: rddata <= 028;
      0956: rddata <= 012;
      0957: rddata <= 000;
      0958: rddata <= 024;
      0959: rddata <= 000;
      0960: rddata <= 003;
      0961: rddata <= 051;
      0962: rddata <= 102;
      0963: rddata <= 099;
      0964: rddata <= 102;
      0965: rddata <= 006;
      0966: rddata <= 006;
      0967: rddata <= 099;
      0968: rddata <= 051;
      0969: rddata <= 012;
      0970: rddata <= 051;
      0971: rddata <= 054;
      0972: rddata <= 102;
      0973: rddata <= 099;
      0974: rddata <= 115;
      0975: rddata <= 099;
      0976: rddata <= 006;
      0977: rddata <= 123;
      0978: rddata <= 102;
      0979: rddata <= 051;
      0980: rddata <= 012;
      0981: rddata <= 051;
      0982: rddata <= 051;
      0983: rddata <= 054;
      0984: rddata <= 051;
      0985: rddata <= 012;
      0986: rddata <= 070;
      0987: rddata <= 012;
      0988: rddata <= 048;
      0989: rddata <= 048;
      0990: rddata <= 000;
      0991: rddata <= 000;
      0992: rddata <= 000;
      0993: rddata <= 051;
      0994: rddata <= 102;
      0995: rddata <= 003;
      0996: rddata <= 051;
      0997: rddata <= 003;
      0998: rddata <= 006;
      0999: rddata <= 051;
      1000: rddata <= 102;
      1001: rddata <= 024;
      1002: rddata <= 048;
      1003: rddata <= 054;
      1004: rddata <= 024;
      1005: rddata <= 107;
      1006: rddata <= 051;
      1007: rddata <= 051;
      1008: rddata <= 102;
      1009: rddata <= 051;
      1010: rddata <= 006;
      1011: rddata <= 024;
      1012: rddata <= 006;
      1013: rddata <= 051;
      1014: rddata <= 051;
      1015: rddata <= 107;
      1016: rddata <= 028;
      1017: rddata <= 102;
      1018: rddata <= 006;
      1019: rddata <= 012;
      1020: rddata <= 024;
      1021: rddata <= 012;
      1022: rddata <= 000;
      1023: rddata <= 099;
      1024: rddata <= 000;
      1025: rddata <= 000;
      1026: rddata <= 195;
      1027: rddata <= 028;
      1028: rddata <= 008;
      1029: rddata <= 024;
      1030: rddata <= 024;
      1031: rddata <= 000;
      1032: rddata <= 000;
      1033: rddata <= 034;
      1034: rddata <= 034;
      1035: rddata <= 051;
      1036: rddata <= 024;
      1037: rddata <= 000;
      1038: rddata <= 231;
      1039: rddata <= 219;
      1040: rddata <= 096;
      1041: rddata <= 003;
      1042: rddata <= 060;
      1043: rddata <= 102;
      1044: rddata <= 216;
      1045: rddata <= 048;
      1046: rddata <= 127;
      1047: rddata <= 060;
      1048: rddata <= 024;
      1049: rddata <= 060;
      1050: rddata <= 000;
      1051: rddata <= 000;
      1052: rddata <= 000;
      1053: rddata <= 000;
      1054: rddata <= 127;
      1055: rddata <= 008;
      1056: rddata <= 000;
      1057: rddata <= 012;
      1058: rddata <= 000;
      1059: rddata <= 054;
      1060: rddata <= 031;
      1061: rddata <= 051;
      1062: rddata <= 059;
      1063: rddata <= 000;
      1064: rddata <= 024;
      1065: rddata <= 012;
      1066: rddata <= 000;
      1067: rddata <= 000;
      1068: rddata <= 028;
      1069: rddata <= 000;
      1070: rddata <= 028;
      1071: rddata <= 003;
      1072: rddata <= 099;
      1073: rddata <= 012;
      1074: rddata <= 051;
      1075: rddata <= 051;
      1076: rddata <= 048;
      1077: rddata <= 051;
      1078: rddata <= 051;
      1079: rddata <= 012;
      1080: rddata <= 051;
      1081: rddata <= 012;
      1082: rddata <= 028;
      1083: rddata <= 028;
      1084: rddata <= 024;
      1085: rddata <= 000;
      1086: rddata <= 012;
      1087: rddata <= 012;
      1088: rddata <= 003;
      1089: rddata <= 051;
      1090: rddata <= 102;
      1091: rddata <= 102;
      1092: rddata <= 054;
      1093: rddata <= 070;
      1094: rddata <= 006;
      1095: rddata <= 102;
      1096: rddata <= 051;
      1097: rddata <= 012;
      1098: rddata <= 051;
      1099: rddata <= 102;
      1100: rddata <= 102;
      1101: rddata <= 099;
      1102: rddata <= 099;
      1103: rddata <= 054;
      1104: rddata <= 006;
      1105: rddata <= 062;
      1106: rddata <= 102;
      1107: rddata <= 051;
      1108: rddata <= 012;
      1109: rddata <= 051;
      1110: rddata <= 030;
      1111: rddata <= 054;
      1112: rddata <= 051;
      1113: rddata <= 012;
      1114: rddata <= 099;
      1115: rddata <= 012;
      1116: rddata <= 096;
      1117: rddata <= 048;
      1118: rddata <= 000;
      1119: rddata <= 000;
      1120: rddata <= 000;
      1121: rddata <= 051;
      1122: rddata <= 102;
      1123: rddata <= 051;
      1124: rddata <= 051;
      1125: rddata <= 051;
      1126: rddata <= 006;
      1127: rddata <= 062;
      1128: rddata <= 102;
      1129: rddata <= 024;
      1130: rddata <= 048;
      1131: rddata <= 102;
      1132: rddata <= 024;
      1133: rddata <= 107;
      1134: rddata <= 051;
      1135: rddata <= 051;
      1136: rddata <= 102;
      1137: rddata <= 051;
      1138: rddata <= 006;
      1139: rddata <= 051;
      1140: rddata <= 054;
      1141: rddata <= 051;
      1142: rddata <= 030;
      1143: rddata <= 054;
      1144: rddata <= 054;
      1145: rddata <= 060;
      1146: rddata <= 035;
      1147: rddata <= 012;
      1148: rddata <= 024;
      1149: rddata <= 012;
      1150: rddata <= 000;
      1151: rddata <= 127;
      1152: rddata <= 000;
      1153: rddata <= 255;
      1154: rddata <= 126;
      1155: rddata <= 008;
      1156: rddata <= 000;
      1157: rddata <= 126;
      1158: rddata <= 126;
      1159: rddata <= 000;
      1160: rddata <= 000;
      1161: rddata <= 028;
      1162: rddata <= 028;
      1163: rddata <= 030;
      1164: rddata <= 024;
      1165: rddata <= 000;
      1166: rddata <= 103;
      1167: rddata <= 024;
      1168: rddata <= 064;
      1169: rddata <= 001;
      1170: rddata <= 024;
      1171: rddata <= 102;
      1172: rddata <= 216;
      1173: rddata <= 099;
      1174: rddata <= 127;
      1175: rddata <= 024;
      1176: rddata <= 024;
      1177: rddata <= 024;
      1178: rddata <= 000;
      1179: rddata <= 000;
      1180: rddata <= 000;
      1181: rddata <= 000;
      1182: rddata <= 127;
      1183: rddata <= 008;
      1184: rddata <= 000;
      1185: rddata <= 012;
      1186: rddata <= 000;
      1187: rddata <= 054;
      1188: rddata <= 012;
      1189: rddata <= 049;
      1190: rddata <= 110;
      1191: rddata <= 000;
      1192: rddata <= 048;
      1193: rddata <= 006;
      1194: rddata <= 000;
      1195: rddata <= 000;
      1196: rddata <= 028;
      1197: rddata <= 000;
      1198: rddata <= 028;
      1199: rddata <= 001;
      1200: rddata <= 062;
      1201: rddata <= 063;
      1202: rddata <= 063;
      1203: rddata <= 030;
      1204: rddata <= 120;
      1205: rddata <= 030;
      1206: rddata <= 030;
      1207: rddata <= 012;
      1208: rddata <= 030;
      1209: rddata <= 014;
      1210: rddata <= 000;
      1211: rddata <= 024;
      1212: rddata <= 048;
      1213: rddata <= 000;
      1214: rddata <= 006;
      1215: rddata <= 012;
      1216: rddata <= 062;
      1217: rddata <= 051;
      1218: rddata <= 063;
      1219: rddata <= 060;
      1220: rddata <= 031;
      1221: rddata <= 127;
      1222: rddata <= 015;
      1223: rddata <= 124;
      1224: rddata <= 051;
      1225: rddata <= 030;
      1226: rddata <= 030;
      1227: rddata <= 103;
      1228: rddata <= 127;
      1229: rddata <= 099;
      1230: rddata <= 099;
      1231: rddata <= 028;
      1232: rddata <= 015;
      1233: rddata <= 048;
      1234: rddata <= 103;
      1235: rddata <= 030;
      1236: rddata <= 030;
      1237: rddata <= 030;
      1238: rddata <= 012;
      1239: rddata <= 054;
      1240: rddata <= 051;
      1241: rddata <= 030;
      1242: rddata <= 127;
      1243: rddata <= 060;
      1244: rddata <= 064;
      1245: rddata <= 060;
      1246: rddata <= 000;
      1247: rddata <= 000;
      1248: rddata <= 000;
      1249: rddata <= 110;
      1250: rddata <= 059;
      1251: rddata <= 030;
      1252: rddata <= 110;
      1253: rddata <= 030;
      1254: rddata <= 015;
      1255: rddata <= 048;
      1256: rddata <= 103;
      1257: rddata <= 126;
      1258: rddata <= 051;
      1259: rddata <= 103;
      1260: rddata <= 126;
      1261: rddata <= 099;
      1262: rddata <= 051;
      1263: rddata <= 030;
      1264: rddata <= 062;
      1265: rddata <= 062;
      1266: rddata <= 015;
      1267: rddata <= 030;
      1268: rddata <= 028;
      1269: rddata <= 110;
      1270: rddata <= 012;
      1271: rddata <= 054;
      1272: rddata <= 099;
      1273: rddata <= 048;
      1274: rddata <= 063;
      1275: rddata <= 056;
      1276: rddata <= 024;
      1277: rddata <= 007;
      1278: rddata <= 000;
      1279: rddata <= 000;
      1280: rddata <= 000;
      1281: rddata <= 000;
      1282: rddata <= 000;
      1283: rddata <= 000;
      1284: rddata <= 000;
      1285: rddata <= 000;
      1286: rddata <= 000;
      1287: rddata <= 000;
      1288: rddata <= 000;
      1289: rddata <= 000;
      1290: rddata <= 000;
      1291: rddata <= 000;
      1292: rddata <= 000;
      1293: rddata <= 000;
      1294: rddata <= 003;
      1295: rddata <= 000;
      1296: rddata <= 000;
      1297: rddata <= 000;
      1298: rddata <= 000;
      1299: rddata <= 000;
      1300: rddata <= 000;
      1301: rddata <= 126;
      1302: rddata <= 000;
      1303: rddata <= 126;
      1304: rddata <= 000;
      1305: rddata <= 000;
      1306: rddata <= 000;
      1307: rddata <= 000;
      1308: rddata <= 000;
      1309: rddata <= 000;
      1310: rddata <= 000;
      1311: rddata <= 000;
      1312: rddata <= 000;
      1313: rddata <= 000;
      1314: rddata <= 000;
      1315: rddata <= 000;
      1316: rddata <= 012;
      1317: rddata <= 000;
      1318: rddata <= 000;
      1319: rddata <= 000;
      1320: rddata <= 000;
      1321: rddata <= 000;
      1322: rddata <= 000;
      1323: rddata <= 000;
      1324: rddata <= 006;
      1325: rddata <= 000;
      1326: rddata <= 000;
      1327: rddata <= 000;
      1328: rddata <= 000;
      1329: rddata <= 000;
      1330: rddata <= 000;
      1331: rddata <= 000;
      1332: rddata <= 000;
      1333: rddata <= 000;
      1334: rddata <= 000;
      1335: rddata <= 000;
      1336: rddata <= 000;
      1337: rddata <= 000;
      1338: rddata <= 000;
      1339: rddata <= 012;
      1340: rddata <= 000;
      1341: rddata <= 000;
      1342: rddata <= 000;
      1343: rddata <= 000;
      1344: rddata <= 000;
      1345: rddata <= 000;
      1346: rddata <= 000;
      1347: rddata <= 000;
      1348: rddata <= 000;
      1349: rddata <= 000;
      1350: rddata <= 000;
      1351: rddata <= 000;
      1352: rddata <= 000;
      1353: rddata <= 000;
      1354: rddata <= 000;
      1355: rddata <= 000;
      1356: rddata <= 000;
      1357: rddata <= 000;
      1358: rddata <= 000;
      1359: rddata <= 000;
      1360: rddata <= 000;
      1361: rddata <= 120;
      1362: rddata <= 000;
      1363: rddata <= 000;
      1364: rddata <= 000;
      1365: rddata <= 000;
      1366: rddata <= 000;
      1367: rddata <= 000;
      1368: rddata <= 000;
      1369: rddata <= 000;
      1370: rddata <= 000;
      1371: rddata <= 000;
      1372: rddata <= 000;
      1373: rddata <= 000;
      1374: rddata <= 000;
      1375: rddata <= 255;
      1376: rddata <= 000;
      1377: rddata <= 000;
      1378: rddata <= 000;
      1379: rddata <= 000;
      1380: rddata <= 000;
      1381: rddata <= 000;
      1382: rddata <= 000;
      1383: rddata <= 051;
      1384: rddata <= 000;
      1385: rddata <= 000;
      1386: rddata <= 051;
      1387: rddata <= 000;
      1388: rddata <= 000;
      1389: rddata <= 000;
      1390: rddata <= 000;
      1391: rddata <= 000;
      1392: rddata <= 006;
      1393: rddata <= 048;
      1394: rddata <= 000;
      1395: rddata <= 000;
      1396: rddata <= 000;
      1397: rddata <= 000;
      1398: rddata <= 000;
      1399: rddata <= 000;
      1400: rddata <= 000;
      1401: rddata <= 024;
      1402: rddata <= 000;
      1403: rddata <= 000;
      1404: rddata <= 000;
      1405: rddata <= 000;
      1406: rddata <= 000;
      1407: rddata <= 000;
      1408: rddata <= 000;
      1409: rddata <= 000;
      1410: rddata <= 000;
      1411: rddata <= 000;
      1412: rddata <= 000;
      1413: rddata <= 000;
      1414: rddata <= 000;
      1415: rddata <= 000;
      1416: rddata <= 000;
      1417: rddata <= 000;
      1418: rddata <= 000;
      1419: rddata <= 000;
      1420: rddata <= 000;
      1421: rddata <= 000;
      1422: rddata <= 000;
      1423: rddata <= 000;
      1424: rddata <= 000;
      1425: rddata <= 000;
      1426: rddata <= 000;
      1427: rddata <= 000;
      1428: rddata <= 000;
      1429: rddata <= 000;
      1430: rddata <= 000;
      1431: rddata <= 000;
      1432: rddata <= 000;
      1433: rddata <= 000;
      1434: rddata <= 000;
      1435: rddata <= 000;
      1436: rddata <= 000;
      1437: rddata <= 000;
      1438: rddata <= 000;
      1439: rddata <= 000;
      1440: rddata <= 000;
      1441: rddata <= 000;
      1442: rddata <= 000;
      1443: rddata <= 000;
      1444: rddata <= 000;
      1445: rddata <= 000;
      1446: rddata <= 000;
      1447: rddata <= 000;
      1448: rddata <= 000;
      1449: rddata <= 000;
      1450: rddata <= 000;
      1451: rddata <= 000;
      1452: rddata <= 000;
      1453: rddata <= 000;
      1454: rddata <= 000;
      1455: rddata <= 000;
      1456: rddata <= 000;
      1457: rddata <= 000;
      1458: rddata <= 000;
      1459: rddata <= 000;
      1460: rddata <= 000;
      1461: rddata <= 000;
      1462: rddata <= 000;
      1463: rddata <= 000;
      1464: rddata <= 000;
      1465: rddata <= 000;
      1466: rddata <= 000;
      1467: rddata <= 000;
      1468: rddata <= 000;
      1469: rddata <= 000;
      1470: rddata <= 000;
      1471: rddata <= 000;
      1472: rddata <= 000;
      1473: rddata <= 000;
      1474: rddata <= 000;
      1475: rddata <= 000;
      1476: rddata <= 000;
      1477: rddata <= 000;
      1478: rddata <= 000;
      1479: rddata <= 000;
      1480: rddata <= 000;
      1481: rddata <= 000;
      1482: rddata <= 000;
      1483: rddata <= 000;
      1484: rddata <= 000;
      1485: rddata <= 000;
      1486: rddata <= 000;
      1487: rddata <= 000;
      1488: rddata <= 000;
      1489: rddata <= 000;
      1490: rddata <= 000;
      1491: rddata <= 000;
      1492: rddata <= 000;
      1493: rddata <= 000;
      1494: rddata <= 000;
      1495: rddata <= 000;
      1496: rddata <= 000;
      1497: rddata <= 000;
      1498: rddata <= 000;
      1499: rddata <= 000;
      1500: rddata <= 000;
      1501: rddata <= 000;
      1502: rddata <= 000;
      1503: rddata <= 000;
      1504: rddata <= 000;
      1505: rddata <= 000;
      1506: rddata <= 000;
      1507: rddata <= 000;
      1508: rddata <= 000;
      1509: rddata <= 000;
      1510: rddata <= 000;
      1511: rddata <= 030;
      1512: rddata <= 000;
      1513: rddata <= 000;
      1514: rddata <= 030;
      1515: rddata <= 000;
      1516: rddata <= 000;
      1517: rddata <= 000;
      1518: rddata <= 000;
      1519: rddata <= 000;
      1520: rddata <= 015;
      1521: rddata <= 120;
      1522: rddata <= 000;
      1523: rddata <= 000;
      1524: rddata <= 000;
      1525: rddata <= 000;
      1526: rddata <= 000;
      1527: rddata <= 000;
      1528: rddata <= 000;
      1529: rddata <= 015;
      1530: rddata <= 000;
      1531: rddata <= 000;
      1532: rddata <= 000;
      1533: rddata <= 000;
      1534: rddata <= 000;
      1535: rddata <= 000;
    endcase

  if (!nRST)
    rddata <= 8'd000;
end

endmodule
